/* Copyright (C) 2025 KEELFW
*
* This library is free software; you can redistribute it and/or
* modify it under the terms of the GNU Lesser General Public
* License as published by the Free Software Foundation; either
* version 2.1 of the License, or (at your option) any later version.
*
* This library is distributed in the hope that it will be useful,
* but WITHOUT ANY WARRANTY; without even the implied warranty of
* MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the GNU
* Lesser General Public License for more details.
*
* You should have received a copy of the GNU Lesser General Public
* License along with this library; if not, write to the Free Software
* Foundation, Inc., 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301  USA
*
* See LICENSE file for full license details.
*
* This code was automatically generated by:
*   axi4lite_reg_generator v1.3.2
*
*/

// Data Size = 32
// Write Strobe Size = 4

module example #(
  parameter ADDRESS_W = 32,
  parameter ADDRESS_APERTURE = 8,
  parameter REGISTER_INPUTS = 0
)(
  input  wire                         REGS_ACLK,
  input  wire                         REGS_ARESETN,
  // Registers
  input wire [31:0] R_Test_Register_I,
  output wire [31:0] R_Scratch_Register_O,
  output reg R_Scratch_Register_O_upd,
  input wire [14:0] R_Register_with_Fields_I,
  output wire [14:0] R_Register_with_Fields_O,
  output reg R_Register_with_Fields_O_upd,
    
  // Write Address Channel
  input  wire                        REGS_AWVALID,
  output reg                         REGS_AWREADY,
  input  wire [ADDRESS_W-1:0]        REGS_AWADDR,
  input  wire [2:0]                  REGS_AWPROT,
  // Write Data Channel
  input  wire                        REGS_WVALID,
  output wire                        REGS_WREADY,
  input  wire [31:0]                 REGS_WDATA,
  input  wire [3:0]                  REGS_WSTRB,
  // Write Response Channel
  output reg                         REGS_BVALID,
  input  wire                        REGS_BREADY,
  output reg  [1:0]                  REGS_BRESP,
  // Read Address Channel
  input  wire                        REGS_ARVALID,
  output reg                         REGS_ARREADY,
  input  wire [ADDRESS_W-1:0]        REGS_ARADDR,
  input  wire [2:0]                  REGS_ARPROT,
  // Read Data Channel
  output wire                        REGS_RVALID,
  input  wire                        REGS_RREADY,
  output reg  [31:0]                 REGS_RDATA,
  output reg  [1:0]                  REGS_RRESP
);

localparam [1:0] AXI_RESP_OKAY   = 2'b00;
localparam [1:0] AXI_RESP_EXOKAY = 2'b01;
localparam [1:0] AXI_RESP_SLVERR = 2'b10;
localparam [1:0] AXI_RESP_DECERR = 2'b11;

// Register signal declarations
reg [31:0] REG_Test_Register_R;

reg [31:0] REG_Scratch_Register_R;
reg [31:0] REG_Scratch_Register_W;

reg [14:0] REG_Register_with_Fields_R;
reg [14:0] REG_Register_with_Fields_W;



// Internal AXI support signals
// Write state machine states
localparam [1:0] W_STATE_RST = 2'b00;
localparam [1:0] W_STATE_WAIT4ADDR = 2'b01;
localparam [1:0] W_STATE_WAIT4DATA = 2'b10;
localparam [1:0] W_STATE_WAIT4RESP = 2'b11;

// Read state machine states
localparam [1:0] R_STATE_RST = 2'b00;
localparam [1:0] R_STATE_WAIT4ADDR = 2'b01;
localparam [1:0] R_STATE_WAITREG = 2'b10;
localparam [1:0] R_STATE_WAIT4DATA = 2'b11;

reg [1:0] state_w;
reg [1:0] state_r;

reg [ADDRESS_APERTURE-1:0] address_wr;
reg [ADDRESS_APERTURE-1:0] address_rd;

reg w_ready;
reg r_valid;

reg [31:0] rd_mux;
reg [1:0] rd_resp;

// Handle inputs

always @* begin
REG_Scratch_Register_R <= REG_Scratch_Register_W;

end

generate
  if (REGISTER_INPUTS > 0) begin : reg_inputs_g
    always @(posedge REGS_ACLK) begin
      REG_Test_Register_R <= R_Test_Register_I; 
      REG_Register_with_Fields_R <= R_Register_with_Fields_I; 
      
    end
  end else begin : con_inputs_g
    always @* begin
      REG_Test_Register_R <= R_Test_Register_I;
      REG_Register_with_Fields_R <= R_Register_with_Fields_I;
      
    end
  end
endgenerate

// Connect outputs
assign R_Scratch_Register_O = REG_Scratch_Register_W;
assign R_Register_with_Fields_O = REG_Register_with_Fields_W;

// Connect AXI-Lite ready/valid control signals
assign REGS_WREADY = w_ready;
assign REGS_RVALID = r_valid;

// Write FSM
always @(posedge REGS_ACLK) begin
  if (!REGS_ARESETN) begin
    state_w <= W_STATE_RST;
    REGS_AWREADY <= 0;
    w_ready <= 0;
    REGS_BVALID <= 0;
  end
  else begin
    case (state_w)
      W_STATE_RST: begin
        state_w <= W_STATE_WAIT4ADDR;
        REGS_AWREADY <= 1;
      end
      W_STATE_WAIT4ADDR: begin
        if (REGS_AWVALID) begin
          state_w <= W_STATE_WAIT4DATA;
          REGS_AWREADY <= 0;
          w_ready <= 1;
          address_wr <= REGS_AWADDR[ADDRESS_APERTURE-1:0];
        end
      end
      W_STATE_WAIT4DATA: begin
        if (REGS_WVALID) begin
          state_w <= W_STATE_WAIT4RESP;
          w_ready <= 0;
          REGS_BVALID <= 1;
        end
      end
      W_STATE_WAIT4RESP: begin
        if (REGS_BREADY) begin
          state_w <= W_STATE_WAIT4ADDR;
          REGS_BVALID <= 0;
          REGS_AWREADY <= 1;
        end
      end
      default: begin
        state_w <= W_STATE_RST;
      end
    endcase
  end
end

// Read FSM
always @(posedge REGS_ACLK) begin
  if (!REGS_ARESETN) begin
    state_r <= R_STATE_RST;
    REGS_ARREADY <= 0;
    r_valid <= 0;
  end
  else begin
    case (state_r)
      R_STATE_RST: begin
        state_r <= R_STATE_WAIT4ADDR;
        REGS_ARREADY <= 1;
      end
      R_STATE_WAIT4ADDR: begin
        if (REGS_ARVALID) begin
          state_r <= R_STATE_WAITREG;
          REGS_ARREADY <= 0;
          address_rd <= REGS_ARADDR[ADDRESS_APERTURE-1:0];
        end
      end
      R_STATE_WAITREG: begin
        state_r <= R_STATE_WAIT4DATA;
        r_valid <= 1;
      end
      R_STATE_WAIT4DATA: begin
        if (REGS_RREADY == 1) begin
          state_r <= R_STATE_WAIT4ADDR;
          r_valid <= 0;
          REGS_ARREADY <= 1;
        end
      end
      default: begin
        state_r <= R_STATE_RST;
      end
    endcase
  end
end

// Write process
always @(posedge REGS_ACLK) begin
  if (!REGS_ARESETN) begin
    REG_Scratch_Register_W <= 32'b00000000000000000000000000000000;
    R_Scratch_Register_O_upd <= 0;
    REG_Register_with_Fields_W <= 15'b011111111110000;
    R_Register_with_Fields_O_upd <= 0;
  end
  else begin
    R_Scratch_Register_O_upd <= 0;
    R_Register_with_Fields_O_upd <= 0;
    if (REGS_WVALID && w_ready) begin
      if (address_wr == 4) begin
        R_Scratch_Register_O_upd <= 1;
        REGS_BRESP <= AXI_RESP_OKAY;
        if (REGS_WSTRB[0] == 1) begin
          REG_Scratch_Register_W[7:0] <= REGS_WDATA[7:0];
        end
        if (REGS_WSTRB[1] == 1) begin
          REG_Scratch_Register_W[15:8] <= REGS_WDATA[15:8];
        end
        if (REGS_WSTRB[2] == 1) begin
          REG_Scratch_Register_W[23:16] <= REGS_WDATA[23:16];
        end
        if (REGS_WSTRB[3] == 1) begin
          REG_Scratch_Register_W[31:24] <= REGS_WDATA[31:24];
        end
      end else if (address_wr == 64) begin
        R_Register_with_Fields_O_upd <= 1;
        REGS_BRESP <= AXI_RESP_OKAY;
        if (REGS_WSTRB[0] == 1) begin
          REG_Register_with_Fields_W[7:0] <= REGS_WDATA[7:0];
        end
        if (REGS_WSTRB[1] == 1) begin
          REG_Register_with_Fields_W[14:8] <= REGS_WDATA[14:8];
        end
      end else begin
        REGS_BRESP <= AXI_RESP_SLVERR;
      end
    end
  end
end

always @* begin
  case (address_rd)
    0: begin
      
      rd_mux = REG_Test_Register_R;
      
      rd_resp = AXI_RESP_OKAY;
    end
    4: begin
      
      rd_mux = REG_Scratch_Register_R;
      
      rd_resp = AXI_RESP_OKAY;
    end
    64: begin
      
      rd_mux = { {17{1'b0}}, REG_Register_with_Fields_R };
      
      rd_resp = AXI_RESP_OKAY;
    end
    
    default: begin
      rd_mux = 0;
      rd_resp = AXI_RESP_SLVERR;
    end
  endcase
end

// Read process
always @(posedge REGS_ACLK) begin
  if (!REGS_ARESETN) begin
  end else begin
    if (state_r == R_STATE_WAITREG) begin
      REGS_RDATA <= rd_mux;
      REGS_RRESP <= rd_resp;
    end
  end
end

endmodule

// SHA-256: ac28d60f95e62d4c9750d35a6cbfc8c07f24e80d843e2982a6bbfe82f1cba6c1