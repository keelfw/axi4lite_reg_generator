/* Copyright (C) 2025 KEELFW
*
* This library is free software; you can redistribute it and/or
* modify it under the terms of the GNU Lesser General Public
* License as published by the Free Software Foundation; either
* version 2.1 of the License, or (at your option) any later version.
*
* This library is distributed in the hope that it will be useful,
* but WITHOUT ANY WARRANTY; without even the implied warranty of
* MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the GNU
* Lesser General Public License for more details.
*
* You should have received a copy of the GNU Lesser General Public
* License along with this library; if not, write to the Free Software
* Foundation, Inc., 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301  USA
*
* See LICENSE file for full license details.
*
* This code was automatically generated by:
*   axi4lite_reg_generator v1.4.0
*
*/

// Data Size = 32
// Write Strobe Size = 4

module example #(
  parameter ADDRESS_W = 32,
  parameter ADDRESS_APERTURE = 8,
  parameter REGISTER_INPUTS = 0
)(
  input  logic                        regs_aclk,
  input  logic                        regs_aresetn,
  // Registers
  input logic [31:0] R_Test_Register_I,
  output logic [31:0] R_Scratch_Register_O,
  output logic R_Scratch_Register_O_upd,
  input logic [14:0] R_Register_with_Fields_I,
  output logic [14:0] R_Register_with_Fields_O,
  output logic R_Register_with_Fields_O_upd,
    
  // Write Address Channel
  input  logic                        regs_awvalid,
  output logic                        regs_awready,
  input  logic [ADDRESS_W-1:0]        regs_awaddr,
  input  logic [2:0]                  regs_awprot,
  // Write Data Channel
  input  logic                        regs_wvalid,
  output logic                        regs_wready,
  input  logic [31:0]                 regs_wdata,
  input  logic [3:0]                  regs_wstrb,
  // Write Response Channel
  output logic                        regs_bvalid,
  input  logic                        regs_bready,
  output logic  [1:0]                 regs_bresp,
  // Read Address Channel
  input  logic                        regs_arvalid,
  output logic                        regs_arready,
  input  logic [ADDRESS_W-1:0]        regs_araddr,
  input  logic [2:0]                  regs_arprot,
  // Read Data Channel
  output logic                        regs_rvalid,
  input  logic                        regs_rready,
  output logic  [31:0]                regs_rdata,
  output logic  [1:0]                 regs_rresp
);

// AXI Response Constants
localparam [1:0] AXI_RESP_OKAY   = 2'b00;
localparam [1:0] AXI_RESP_EXOKAY = 2'b01;
localparam [1:0] AXI_RESP_SLVERR = 2'b10;
localparam [1:0] AXI_RESP_DECERR = 2'b11;

// Register addresses
localparam [ADDRESS_APERTURE-1:0] REG_Test_Register_ADDR = 0;
localparam [ADDRESS_APERTURE-1:0] REG_Scratch_Register_ADDR = 4;
localparam [ADDRESS_APERTURE-1:0] REG_Register_with_Fields_ADDR = 64;


// Register signal declarations
logic [31:0] REG_Test_Register_R;

logic [31:0] REG_Scratch_Register_R;
logic [31:0] REG_Scratch_Register_W;

logic [14:0] REG_Register_with_Fields_R;
logic [14:0] REG_Register_with_Fields_W;



// Internal AXI support signals
// Write state machine states
typedef enum logic [1:0] {
    W_STATE_RST,
    W_STATE_WAIT4ADDR,
    W_STATE_WAIT4DATA,
    W_STATE_WAIT4RESP
} write_state_t;

// Read state machine states
typedef enum logic [1:0] {
    R_STATE_RST,
    R_STATE_WAIT4ADDR,
    R_STATE_WAITREG,
    R_STATE_WAIT4DATA
} read_state_t;

write_state_t state_w;
read_state_t state_r;

logic [ADDRESS_APERTURE-1:0] address_wr;
logic [ADDRESS_APERTURE-1:0] address_rd;

logic w_ready;
logic r_valid;

logic [31:0] rd_mux;
logic [1:0] rd_resp;

// Handle inputs

always_comb begin
REG_Scratch_Register_R = REG_Scratch_Register_W;

end

generate
  if (REGISTER_INPUTS > 0) begin : reg_inputs_g
    always_ff @(posedge regs_aclk) begin
      REG_Test_Register_R <= R_Test_Register_I; 
      REG_Register_with_Fields_R <= R_Register_with_Fields_I; 
      
    end
  end else begin : con_inputs_g
    always_comb begin
      REG_Test_Register_R = R_Test_Register_I;
      REG_Register_with_Fields_R = R_Register_with_Fields_I;
      
    end
  end
endgenerate

// Connect outputs
assign R_Scratch_Register_O = REG_Scratch_Register_W;
assign R_Register_with_Fields_O = REG_Register_with_Fields_W;

// Connect AXI-Lite ready/valid control signals
assign regs_wready = w_ready;
assign regs_rvalid = r_valid;

// Write FSM
always_ff @(posedge regs_aclk) begin
  if (!regs_aresetn) begin
    state_w <= W_STATE_RST;
    regs_awready <= '0;
    w_ready <= '0;
    regs_bvalid <= '0;
  end
  else begin
    case (state_w)
      W_STATE_RST: begin
        state_w <= W_STATE_WAIT4ADDR;
        regs_awready <= '1;
      end
      W_STATE_WAIT4ADDR: begin
        if (regs_awvalid) begin
          state_w <= W_STATE_WAIT4DATA;
          regs_awready <= '0;
          w_ready <= '1;
          address_wr <= regs_awaddr[ADDRESS_APERTURE-1:0];
        end
      end
      W_STATE_WAIT4DATA: begin
        if (regs_wvalid) begin
          state_w <= W_STATE_WAIT4RESP;
          w_ready <= '0;
          regs_bvalid <= '1;
        end
      end
      W_STATE_WAIT4RESP: begin
        if (regs_bready) begin
          state_w <= W_STATE_WAIT4ADDR;
          regs_bvalid <= '0;
          regs_awready <= '1;
        end
      end
      default: begin
        state_w <= W_STATE_RST;
      end
    endcase
  end
end

// Read FSM
always_ff @(posedge regs_aclk) begin
  if (!regs_aresetn) begin
    state_r <= R_STATE_RST;
    regs_arready <= '0;
    r_valid <= '0;
  end
  else begin
    case (state_r)
      R_STATE_RST: begin
        state_r <= R_STATE_WAIT4ADDR;
        regs_arready <= '1;
      end
      R_STATE_WAIT4ADDR: begin
        if (regs_arvalid) begin
          state_r <= R_STATE_WAITREG;
          regs_arready <= '0;
          address_rd <= regs_araddr[ADDRESS_APERTURE-1:0];
        end
      end
      R_STATE_WAITREG: begin
        state_r <= R_STATE_WAIT4DATA;
        r_valid <= '1;
      end
      R_STATE_WAIT4DATA: begin
        if (regs_rready) begin
          state_r <= R_STATE_WAIT4ADDR;
          r_valid <= '0;
          regs_arready <= '1;
        end
      end
      default: begin
        state_r <= R_STATE_RST;
      end
    endcase
  end
end

// Write process
always_ff @(posedge regs_aclk) begin
  if (!regs_aresetn) begin
    REG_Scratch_Register_W <= 32'b00000000000000000000000000000000;
    R_Scratch_Register_O_upd <= '0;
    REG_Register_with_Fields_W <= 15'b011111111110000;
    R_Register_with_Fields_O_upd <= '0;
  end
  else begin
    R_Scratch_Register_O_upd <= '0;
    R_Register_with_Fields_O_upd <= '0;
    if (regs_wvalid && w_ready) begin
      if (address_wr == REG_Scratch_Register_ADDR) begin
        R_Scratch_Register_O_upd <= '1;
        regs_bresp <= AXI_RESP_OKAY;
        if (regs_wstrb[0]) begin
          REG_Scratch_Register_W[7:0] <= regs_wdata[7:0];
        end
        if (regs_wstrb[1]) begin
          REG_Scratch_Register_W[15:8] <= regs_wdata[15:8];
        end
        if (regs_wstrb[2]) begin
          REG_Scratch_Register_W[23:16] <= regs_wdata[23:16];
        end
        if (regs_wstrb[3]) begin
          REG_Scratch_Register_W[31:24] <= regs_wdata[31:24];
        end
      end else if (address_wr == REG_Register_with_Fields_ADDR) begin
        R_Register_with_Fields_O_upd <= '1;
        regs_bresp <= AXI_RESP_OKAY;
        if (regs_wstrb[0]) begin
          REG_Register_with_Fields_W[7:0] <= regs_wdata[7:0];
        end
        if (regs_wstrb[1]) begin
          REG_Register_with_Fields_W[14:8] <= regs_wdata[14:8];
        end
      end else begin
        regs_bresp <= AXI_RESP_SLVERR;
      end
    end
  end
end

always_comb begin
  case (address_rd)
    REG_Test_Register_ADDR: begin
      
      rd_mux = REG_Test_Register_R;
      
      rd_resp = AXI_RESP_OKAY;
    end
    REG_Scratch_Register_ADDR: begin
      
      rd_mux = REG_Scratch_Register_R;
      
      rd_resp = AXI_RESP_OKAY;
    end
    REG_Register_with_Fields_ADDR: begin
      
      rd_mux = { {17{1'b0}}, REG_Register_with_Fields_R };
      
      rd_resp = AXI_RESP_OKAY;
    end
    
    default: begin
      rd_mux = '0;
      rd_resp = AXI_RESP_SLVERR;
    end
  endcase
end

// Read process
always_ff @(posedge regs_aclk) begin
  if (!regs_aresetn) begin
  end else begin
    if (state_r == R_STATE_WAITREG) begin
      regs_rdata <= rd_mux;
      regs_rresp <= rd_resp;
    end
  end
end

endmodule

// SHA-256: eea38166ca79f39bbd43eeefcf6b40e4db4ba5a54c576d607b75929fe586c8ad