/* Copyright (C) 2025 KEELFW
*
* This library is free software; you can redistribute it and/or
* modify it under the terms of the GNU Lesser General Public
* License as published by the Free Software Foundation; either
* version 2.1 of the License, or (at your option) any later version.
*
* This library is distributed in the hope that it will be useful,
* but WITHOUT ANY WARRANTY; without even the implied warranty of
* MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the GNU
* Lesser General Public License for more details.
*
* You should have received a copy of the GNU Lesser General Public
* License along with this library; if not, write to the Free Software
* Foundation, Inc., 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301  USA
*
* See LICENSE file for full license details.
*
* This code was automatically generated by:
*   axi4lite_reg_generator v{{ id_version }}
*{% if include_username or include_hostname %} generated by: {% if include_username %}{{ id_username }}{% endif %}{% if include_hostname %}@{{ id_hostname }}{% endif %}{% endif %}{% if include_timestamp %} at {{ id_timestamp }}{% endif %}
*/

// Data Size = {{ data_size }}
// Write Strobe Size = {{ strobe_size }}

module {{ entity_name }} #(
  parameter ADDRESS_W = 32,
  parameter ADDRESS_APERTURE = 8,
  parameter REGISTER_INPUTS = 0
)(
  input  logic                        regs_aclk,
  input  logic                        regs_aresetn,
  // Registers
  {% for reg in regs -%}
  {% if reg['reg_type'] == 'ro' or reg['reg_type'] == 'custom' -%}
  input logic [{{ reg['bits']|count_bits - 1 }}:0] R_{{ reg['name'] }}_I,
  {% endif -%}
  {% if reg['reg_type'] == 'rw' or reg['reg_type'] == 'custom' -%}
  output logic [{{ reg['bits']|count_bits - 1 }}:0] R_{{ reg['name'] }}_O,
  {% if reg['use_upd_pulse'] -%}
  output logic R_{{ reg['name'] }}_O_upd,
  {% endif -%}
  {% endif -%}
  {% endfor %}  
  // Write Address Channel
  input  logic                        regs_awvalid,
  output logic                        regs_awready,
  input  logic [ADDRESS_W-1:0]        regs_awaddr,
  input  logic [2:0]                  regs_awprot,
  // Write Data Channel
  input  logic                        regs_wvalid,
  output logic                        regs_wready,
  input  logic [31:0]                 regs_wdata,
  input  logic [3:0]                  regs_wstrb,
  // Write Response Channel
  output logic                        regs_bvalid,
  input  logic                        regs_bready,
  output logic  [1:0]                 regs_bresp,
  // Read Address Channel
  input  logic                        regs_arvalid,
  output logic                        regs_arready,
  input  logic [ADDRESS_W-1:0]        regs_araddr,
  input  logic [2:0]                  regs_arprot,
  // Read Data Channel
  output logic                        regs_rvalid,
  input  logic                        regs_rready,
  output logic  [31:0]                regs_rdata,
  output logic  [1:0]                 regs_rresp
);

// AXI Response Constants
localparam [1:0] AXI_RESP_OKAY   = 2'b00;
localparam [1:0] AXI_RESP_EXOKAY = 2'b01;
localparam [1:0] AXI_RESP_SLVERR = 2'b10;
localparam [1:0] AXI_RESP_DECERR = 2'b11;

// Register addresses
{% for reg in regs -%}
localparam [ADDRESS_APERTURE-1:0] REG_{{ reg['name'] }}_ADDR = {{ reg['addr_offset'] }};
{% endfor %}

// Register signal declarations
{% for reg in regs -%}
logic [{{ reg['bits']|count_bits-1}}:0] REG_{{ reg['name'] }}_R;
{% if reg['reg_type'] == 'rw' or reg['reg_type'] == 'custom' -%}
logic [{{ reg['bits']|count_bits-1 }}:0] REG_{{ reg['name'] }}_W;
{% endif %}
{% endfor %}

// Internal AXI support signals
// Write state machine states
typedef enum logic [1:0] {
    W_STATE_RST,
    W_STATE_WAIT4ADDR,
    W_STATE_WAIT4DATA,
    W_STATE_WAIT4RESP
} write_state_t;

// Read state machine states
typedef enum logic [1:0] {
    R_STATE_RST,
    R_STATE_WAIT4ADDR,
    R_STATE_WAITREG,
    R_STATE_WAIT4DATA
} read_state_t;

write_state_t state_w;
read_state_t state_r;

logic [ADDRESS_APERTURE-1:0] address_wr;
logic [ADDRESS_APERTURE-1:0] address_rd;

logic w_ready;
logic r_valid;

logic [{{ data_size-1 }}:0] rd_mux;
logic [1:0] rd_resp;

// Handle inputs

always_comb begin
{% for reg in regs -%}
{% if reg['reg_type'] == 'rw' -%}
  REG_{{ reg['name'] }}_R = REG_{{ reg['name'] }}_W;
{% endif -%}
{% endfor %}
end

generate
  if (REGISTER_INPUTS > 0) begin : reg_inputs_g
    always_ff @(posedge regs_aclk) begin
      {% for reg in regs -%}
      {% if reg['reg_type'] == 'ro' or reg['reg_type'] == 'custom' -%}
        REG_{{ reg['name'] }}_R <= R_{{ reg['name'] }}_I; 
      {% endif -%}
      {% endfor %}
    end
  end else begin : con_inputs_g
    always_comb begin
      {% for reg in regs -%}
      {% if reg['reg_type'] != 'rw' -%}
        REG_{{ reg['name'] }}_R = R_{{ reg['name'] }}_I;
      {% endif -%}
      {% endfor %}
    end
  end
endgenerate

// Connect outputs
{% for reg in regs -%}
{% if reg['reg_type'] == 'rw' or reg['reg_type'] == 'custom' -%}
  assign R_{{ reg['name'] }}_O = REG_{{ reg['name'] }}_W;
{% endif -%}
{% endfor %}
// Connect AXI-Lite ready/valid control signals
assign regs_wready = w_ready;
assign regs_rvalid = r_valid;

// Write FSM
always_ff @(posedge regs_aclk) begin
  if (!regs_aresetn) begin
    state_w <= W_STATE_RST;
    regs_awready <= '0;
    w_ready <= '0;
    regs_bvalid <= '0;
  end
  else begin
    case (state_w)
      W_STATE_RST: begin
        state_w <= W_STATE_WAIT4ADDR;
        regs_awready <= '1;
      end
      W_STATE_WAIT4ADDR: begin
        if (regs_awvalid) begin
          state_w <= W_STATE_WAIT4DATA;
          regs_awready <= '0;
          w_ready <= '1;
          address_wr <= regs_awaddr[ADDRESS_APERTURE-1:0];
        end
      end
      W_STATE_WAIT4DATA: begin
        if (regs_wvalid) begin
          state_w <= W_STATE_WAIT4RESP;
          w_ready <= '0;
          regs_bvalid <= '1;
        end
      end
      W_STATE_WAIT4RESP: begin
        if (regs_bready) begin
          state_w <= W_STATE_WAIT4ADDR;
          regs_bvalid <= '0;
          regs_awready <= '1;
        end
      end
      default: begin
        state_w <= W_STATE_RST;
      end
    endcase
  end
end

// Read FSM
always_ff @(posedge regs_aclk) begin
  if (!regs_aresetn) begin
    state_r <= R_STATE_RST;
    regs_arready <= '0;
    r_valid <= '0;
  end
  else begin
    case (state_r)
      R_STATE_RST: begin
        state_r <= R_STATE_WAIT4ADDR;
        regs_arready <= '1;
      end
      R_STATE_WAIT4ADDR: begin
        if (regs_arvalid) begin
          state_r <= R_STATE_WAITREG;
          regs_arready <= '0;
          address_rd <= regs_araddr[ADDRESS_APERTURE-1:0];
        end
      end
      R_STATE_WAITREG: begin
        state_r <= R_STATE_WAIT4DATA;
        r_valid <= '1;
      end
      R_STATE_WAIT4DATA: begin
        if (regs_rready) begin
          state_r <= R_STATE_WAIT4ADDR;
          r_valid <= '0;
          regs_arready <= '1;
        end
      end
      default: begin
        state_r <= R_STATE_RST;
      end
    endcase
  end
end

// Write process
always_ff @(posedge regs_aclk) begin
  if (!regs_aresetn) begin
    {%- for reg in regs -%}
    {%- if reg['reg_type'] == 'rw' or reg['reg_type'] == 'custom' %}
    REG_{{ reg['name'] }}_W <= {{ reg|default_val_v }};
    {%- if reg['use_upd_pulse'] %}
    R_{{ reg['name'] }}_O_upd <= '0;
    {%- endif %}
    {%- endif %}
    {%- endfor %}
  end
  else begin
    {%- for reg in regs -%}
    {%- if reg['reg_type'] == 'rw' or reg['reg_type'] == 'custom' %}
    {%- if reg['use_upd_pulse'] %}
    R_{{ reg['name'] }}_O_upd <= '0;
    {%- endif %}
    {%- endif %}
    {%- endfor %}
    if (regs_wvalid && w_ready) begin
      {% for reg in regs -%}
      {% if reg['reg_type'] == 'rw' or reg['reg_type'] == 'custom' -%}
      if (address_wr == REG_{{ reg['name'] }}_ADDR) begin
        {%- if reg['use_upd_pulse'] %}
        R_{{ reg['name'] }}_O_upd <= '1;
        {%- endif %}
        regs_bresp <= AXI_RESP_OKAY;
        {%- for s in range(strobe_size) %}
        {%- if 8*s < reg['bits']|count_bits %}
        if (regs_wstrb[{{s}}]) begin
          REG_{{ reg['name'] }}_W[{{ [reg['bits']|count_bits-1, 8*(s+1)-1]|min }}:{{ 8*s }}] <= regs_wdata[{{ [reg['bits']|count_bits-1, 8*(s+1)-1]|min }}:{{ 8*s }}];
        end
        {%- endif %}
        {%- endfor %}
      end else {% endif -%}{% endfor -%} begin
        regs_bresp <= AXI_RESP_SLVERR;
      end
    end
  end
end

always_comb begin
  case (address_rd)
    {% for reg in regs -%}
    REG_{{ reg['name'] }}_ADDR: begin
      {% if reg['bits']|count_bits < data_size %}
      rd_mux = {{'{ {'}}{{ data_size - reg['bits']|count_bits }}{1'b0{{'}}'}}, REG_{{ reg['name'] }}_R };
      {% else %}
      rd_mux = REG_{{ reg['name'] }}_R;
      {% endif %}
      rd_resp = AXI_RESP_OKAY;
    end
    {% endfor %}
    default: begin
      rd_mux = '0;
      rd_resp = AXI_RESP_SLVERR;
    end
  endcase
end

// Read process
always_ff @(posedge regs_aclk) begin
  if (!regs_aresetn) begin
  end else begin
    if (state_r == R_STATE_WAITREG) begin
      regs_rdata <= rd_mux;
      regs_rresp <= rd_resp;
    end
  end
end

endmodule

